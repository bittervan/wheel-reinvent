module top (
    output wire led
);

assign led = 1;

endmodule